/******************************************************************
* Description
*	This is an 32-bit arithetic logic unit that can execute the next set of operations:
*		add
*		sub
*		or
*		and
*		nor
* This ALU is written by using behavioral description.
* Version:
*	1.0
* Author:
*	Dr. José Luis Pizano Escalante
* email:
*	luispizano@iteso.mx
* Date:
*	01/03/2014
******************************************************************/
module ALU 
(
	input [3:0] ALUOperation,
	input [31:0] A,
	input [31:0] B,
	input [4:0]shamt, //se agregó debido a que para las operaciones de shift se necesita esta parte de información
	output reg Zero,
	output reg [31:0]ALUResult
);
localparam AND = 4'b0000;
localparam OR  = 4'b0001;
localparam NOR = 4'b0010;
localparam ADD = 4'b0011;
localparam SUB = 4'b0100;

localparam LUI = 4'b0101; //proveniente de alucontrol
localparam Sll = 4'b1111; //proveniente de alucontrol
localparam Srl = 4'b1110;//proveniente de alucontrol


   
   always @ (A or B or ALUOperation)
     begin
		case (ALUOperation)
		  ADD: // add
			ALUResult = A + B;
			
		  SUB:
			ALUResult= A-B;
		  
		  AND:
		  ALUResult= A & B;
			
 		  OR: // or
			ALUResult = A | B;
			
		  NOR: // Nor
			ALUResult = ~(A | B);	
 
		  LUI: //lui agregado 
		   ALUResult = {B[15:0],16'b0000000000000000};	
			
		  Srl: //srl recorrer n bits a la derecha
			ALUResult = B >> shamt;
			
		  Sll: //sll recorrer n bits a la izquierda
			ALUResult = B << shamt;
  
		default:
			ALUResult= 0;
		endcase // case(control)
		Zero = (ALUResult==0) ? 1'b1 : 1'b0;
     end // always @ (A or B or control)
endmodule // ALU